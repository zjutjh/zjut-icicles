LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY CONTROL IS
	PORT(SW0,SW1:IN STD_LOGIC;
		  IN1,IN2,IN3:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		  OU:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		  );
END CONTROL;

ARCHITECTURE one OF CONTROL IS
BEGIN
	PROCESS(SW0,SW1)
	BEGIN
		IF(SW0='0')THEN
			IF(SW1='0')THEN
				OU<=IN1;
			ELSE
				OU<=IN1;
			END IF;
		END IF;
		IF(SW0='1')THEN
			IF(SW1='0')THEN
				OU<=IN2;
			ELSE
				OU<=IN3;
			END IF;
		END IF;
	END PROCESS;
END one;