LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY chose IS
	PORT(keycnt:IN STD_LOGIC;
		  CLK: IN STD_LOGIC;
		  control:OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		  LEDA,LEDB:OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		  );
END chose;

ARCHITECTURE one OF chose IS
	SIGNAL q:STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN
	PROCESS(keycnt)
	BEGIN
		IF(keycnt'EVENT AND keycnt='0')THEN
			IF(q=30)THEN
				q<="00000";
			ELSE
				q<=q+3 after 50ms;
			END IF;
		END IF;
	END PROCESS;
	PROCESS(q)
	BEGIN
		CASE q IS
			WHEN"00000"=>
			control<=X"00029F17";LEDA<="0000110";LEDB<="0111111";
			WHEN"00001"=>
			control<=X"00053E2E";LEDA<="1011011";LEDB<="0111111";
			WHEN"00010"=>
			control<=X"0007DD45";LEDA<="1001111";LEDB<="0111111";
			WHEN"00011"=>
			control<=X"000A7C5C";LEDA<="1100110";LEDB<="0111111";
			WHEN"00100"=>
			control<=X"000D1B71";LEDA<="1101101";LEDB<="0111111";
			WHEN"00101"=>
			control<=X"000FBA8A";LEDA<="1111101";LEDB<="0111111";
			WHEN"00110"=>
			control<=X"001259A1";LEDA<="0000111";LEDB<="0111111";
			WHEN"00111"=>
			control<=X"0014F8B8";LEDA<="1111111";LEDB<="0111111";
			WHEN"01000"=>
			control<=X"001797CF";LEDA<="1101111";LEDB<="0111111";
			WHEN"01001"=>
			control<=X"001A36E6";LEDA<="0111111";LEDB<="0000110";
			WHEN"01010"=>
			control<=X"001CD5FD";LEDA<="0000110";LEDB<="0000110";
			WHEN"01011"=>
			control<=X"001F7514";LEDA<="1011011";LEDB<="0000110";
			WHEN"01100"=>
			control<=X"0022142B";LEDA<="1001111";LEDB<="0000110";
			WHEN"01101"=>
			control<=X"0024B342";LEDA<="1100110";LEDB<="0000110";
			WHEN"01110"=>
			control<=X"00275259";LEDA<="1101101";LEDB<="0000110";
			WHEN"01111"=>
			control<=X"0029F170";LEDA<="1111101";LEDB<="0000110";
			WHEN"10000"=>
			control<=X"002C9087";LEDA<="0000111";LEDB<="0000110";
			WHEN"10001"=>
			control<=X"002F2F9E";LEDA<="1111111";LEDB<="0000110";
			WHEN"10010"=>
			control<=X"0031CEB5";LEDA<="1101111";LEDB<="0000110";
			WHEN"10011"=>
			control<=X"00346DCC";LEDA<="0111111";LEDB<="1011011";
			WHEN"10100"=>
			control<=X"00370CE3";LEDA<="0000110";LEDB<="1011011";
			WHEN"10101"=>
			control<=X"0039ABFA";LEDA<="1011011";LEDB<="1011011";
			WHEN"10110"=>
			control<=X"003C4B11";LEDA<="1001111";LEDB<="1011011";
			WHEN"10111"=>
			control<=X"003EEA28";LEDA<="1100110";LEDB<="1011011";
			WHEN"11000"=>
			control<=X"0041893F";LEDA<="1101101";LEDB<="1011011";
			WHEN"11001"=>
			control<=X"00442856";LEDA<="1111101";LEDB<="1011011";
			WHEN"11010"=>
			control<=X"0046C76D";LEDA<="0000111";LEDB<="1011011";
			WHEN"11011"=>
			control<=X"00496684";LEDA<="1111111";LEDB<="1011011";
			WHEN"11100"=>
			control<=X"004C059B";LEDA<="1101111";LEDB<="1011011";
			WHEN"11101"=>
			control<=X"004EA4B2";LEDA<="0111111";LEDB<="1001111";
			WHEN"11110"=>
			control<=X"005143C9";LEDA<="0000110";LEDB<="1001111";
			WHEN"11111"=>
			control<=X"0053E2E0";LEDA<="1011011";LEDB<="1001111";
			WHEN OTHERS=>
			control<=X"00029F17";LEDA<="0000110";LEDB<="0111111";
		END CASE;
	END PROCESS;
END one;