LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY PHASE_ACC IS
	PORT(clk:IN STD_LOGIC;
		  freqin:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		  romaddr:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		  );
END PHASE_ACC;

ARCHITECTURE  one OF PHASE_ACC IS
		SIGNAL acc:STD_LOGIC_VECTOR(31 DOWNTO 0);
		BEGIN
		PROCESS(clk)
		BEGIN
			IF(clk'EVENT AND clk='1')THEN
				acc<=acc+freqin;
			END IF;
		END PROCESS;
		romaddr<=acc(31 DOWNTO 24);
END one;